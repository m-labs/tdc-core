-------------------------------------------------------------------------------
-- TDC Core / CERN
-------------------------------------------------------------------------------
--
-- unit name: tb_lbc
--
-- author: Sebastien Bourdeauducq, sebastien@milkymist.org
--
-- description: Test bench for leading bit counter
--
-- references: http://www.ohwr.org/projects/tdc-core
--
-------------------------------------------------------------------------------
-- last changes:
-- 2011-08-03 SB Created file
-------------------------------------------------------------------------------

-- Copyright (C) 2011 Sebastien Bourdeauducq

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity tb_lbc is
    generic(
        g_N: positive := 6
    );
end entity;

architecture tb of tb_lbc is

function chr(sl: std_logic) return character is
variable v_c: character;
begin
    case sl is
        when 'U' => v_c:= 'U';
        when 'X' => v_c:= 'X';
        when '0' => v_c:= '0';
        when '1' => v_c:= '1';
        when 'Z' => v_c:= 'Z';
        when 'W' => v_c:= 'W';
        when 'L' => v_c:= 'L';
        when 'H' => v_c:= 'H';
        when '-' => v_c:= '-';
    end case;
return v_c;
end function;

function str(slv: std_logic_vector) return string is
variable result : string (1 to slv'length);
variable r      : integer;
begin
    r := 1;
    for i in slv'range loop
        result(r) := chr(slv(i));
        r := r + 1;
    end loop;
    return result;
end function;

signal clk      : std_logic;
signal polarity : std_logic;
signal d        : std_logic_vector(2**g_N-2 downto 0);
signal count    : std_logic_vector(g_N-1 downto 0);

begin
    dut: entity work.tdc_lbc
        generic map(
            g_N => g_N
        )
        port map(
            clk_i        => clk,
            polarity_i   => polarity,
            d_i          => d,
            count_o      => count
        );
    polarity <= '0';
    process
    variable v_seed1     : positive := 1;
    variable v_seed2     : positive := 2;
    variable v_rand      : real;
    variable v_int_rand  : integer;
    variable v_stim      : std_logic_vector(0 downto 0); 
    begin
        for i in 0 to 2**g_N-1 loop
            -- generate test vector
            for j in 0 to 2**g_N-2 loop
                if j > 2**g_N-2-i then
                    d(j) <= '1';
                elsif j = 2**g_N-2-i then
                    d(j) <= '0';
                else
                    uniform(v_seed1, v_seed2, v_rand);
                    v_int_rand := integer(trunc(v_rand*2.0));
                    v_stim := std_logic_vector(to_unsigned(v_int_rand, v_stim'length));
                    d(j) <= v_stim(0);
                end if;
            end loop;
            -- generate, print and verify output
            clk <= '0';
            wait for 4 ns;
            clk <= '1';
            wait for 4 ns;
            report "Vector:" & str(d) & " Expected:" & integer'image(i) & " Result:" & integer'image(to_integer(unsigned(count)));
            assert i = to_integer(unsigned(count)) severity failure;
        end loop;
        report "Test passed.";
        wait;
    end process;
end architecture;
